// ---********************************************************************------
// Copyright 2020-2030 (c) , Inc. All rights reserved.
// Module Name:   mips_clz.v
// Author     :   tianshuo@firefox.com
// Project Name:  SOC_CBB
// Create Date:   2023-03-26
// Description:
//
// ---********************************************************************------
`ifndef _MIPS_CLZ_V__
`define _MIPS_CLZ_V__

module mips_clz
   #(
    parameter DATA_WIDTH                       = 32,
    parameter DATA_WIDTH_LOG2                  = 5
    )
    (
    input                       [DATA_WIDTH-1:0] data_i,
    output reg               [DATA_WIDTH_LOG2:0] res_o
    );
// -----------------------------------------------------------------------------
// Constant Parameter
// -----------------------------------------------------------------------------

// -----------------------------------------------------------------------------
// Internal Signals Declarations
// -----------------------------------------------------------------------------

// -----------------------------------------------------------------------------
// Main Code
// -----------------------------------------------------------------------------
// ---->TODO
always @(*)
begin
  integer i;
  res_o                      = {1'b1, {DATA_WIDTH_LOG2{1'b0}}};
  for (i = DATA_WIDTH-1; i >= 0; i = i - 1)
  begin
    if (data_i[DATA_WIDTH-1-i] == 1'b1)
      res_o                  = {1'b0, i[DATA_WIDTH_LOG2-1:0]};
  end
end

// -----------------------------------------------------------------------------
// Assertion Declarations
// -----------------------------------------------------------------------------
`ifdef SOC_ASSERT_ON

`endif
endmodule
`endif

// ---********************************************************************------
