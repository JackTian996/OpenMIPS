// ---********************************************************************------
// Copyright 2020-2030 (c) , Inc. All rights reserved.
// Module Name:   LLbit_reg.v
// Author     :   tianshuo@firefox.com
// Project Name:  OPEN_MIPS
// Create Date:   2023-04-09
// Description:
//
// ---********************************************************************------
module llbit_reg
    (
    input                                        clk,
    input                                        rst_n,
    input                                        flush,                        // exception trigger
    input                                        we,
    input                                        llbit_i,
    output reg                                   llbit_o
    );
// -----------------------------------------------------------------------------
// Constant Parameter
// -----------------------------------------------------------------------------

// -----------------------------------------------------------------------------
// Internal Signals Declarations
// -----------------------------------------------------------------------------

// -----------------------------------------------------------------------------
// Main Code
// -----------------------------------------------------------------------------
// ---->TODO
always @(posedge clk or negedge rst_n)
begin : LLBIT_O_PROC
  if (rst_n == `RstEnable)
    llbit_o                  <= {1{1'b0}};
  else if (flush == 1'b1)
    llbit_o                  <= {1{1'b0}};
  else if (we == `WriteEnable)
    llbit_o                  <= llbit_i;
end

// -----------------------------------------------------------------------------
// Assertion Declarations
// -----------------------------------------------------------------------------
`ifdef SOC_ASSERT_ON

`endif
endmodule

// ---********************************************************************------
