// ---********************************************************************------
// Copyright 2020-2030 (c) , Inc. All rights reserved.
// Module Name:   stall_ctrl.v
// Author     :   tianshuo@firefox.com
// Project Name:  OPEN_MIPS
// Create Date:   2023-03-29
// Description:
//
// ---********************************************************************------
module stall_ctrl
    (
    input                                        rst_n,
    input                                        stallreq_from_id,
    input                                        stallreq_from_ex,
    output reg                             [5:0] stall
    );
// -----------------------------------------------------------------------------
// Constant Parameter
// -----------------------------------------------------------------------------

// -----------------------------------------------------------------------------
// Internal Signals Declarations
// -----------------------------------------------------------------------------

// -----------------------------------------------------------------------------
// Main Code
// -----------------------------------------------------------------------------
// ---->TODO

always @(*)
begin : STALL_PROC
  if (rst_n == `RstEnable)
    stall                    = {6{1'b0}};
  else if (stallreq_from_ex == `Stop)
    stall                    = 6'b001111;
  else if (stallreq_from_id == `Stop)
    stall                    = 6'b000111;
  else
    stall                    = {6{1'b0}};
end



// -----------------------------------------------------------------------------
// Assertion Declarations
// -----------------------------------------------------------------------------
`ifdef SOC_ASSERT_ON

`endif
endmodule

// ---********************************************************************------
